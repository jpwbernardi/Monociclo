library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Controle is
  Port(
    bla: in std_logic
  );
end Controle;

architecture cmp of Controle is
begin
end cmp;
