
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.NovosTipos.ALL;

entity tb_mips2 is
end tb_mips2;

architecture cmp of tb_mips2 is
  
  component MIPS is
    Port(
      programa: in VetorWord(0 to 63);
      clk, reset: in std_logic
    );
  end component;
  
signal pro: VetorWord(0 to 63);
signal clock, rst: std_logic;
  
begin
  
  testa: MIPS port map(pro, clock, rst);
  
  --Demonstrando que comando de lw e sw funcionam, j� que n�o fizemos o c�digo do sort
  
  process
  begin
    rst <= '1';
    wait for 2 ns;
    rst <= '0';
   clock <= '0';
    
   pro(0) <= "00000000000000000100000000100000";
   pro(1) <= "00100000000010010000000000001000"; 
   pro(2) <= "10101101000010010000000000000000"; 
  	pro(3) <= "00100001000010000000000000001000"; 
  	pro(4) <= "00100000000010010000000000000010"; 
  	pro(5) <= "10101101000010010000000000000000"; 
  	pro(6) <= "00100001000010000000000000001000"; 
  	pro(7) <= "00100000000010010000000000000111"; 
  	pro(8) <= "10101101000010010000000000000000"; 
  	pro(9) <= "00100001000010000000000000001000";
  	pro(10) <= "00100000000010010000000000001001"; 
  	pro(11) <= "10101101000010010000000000000000";
  	pro(12) <= "00100001000010000000000000001000";
  	pro(13) <= "00100000000010010000000000001000";
  	pro(14) <= "10101101000010010000000000000000";
  	pro(15) <= "00100001000010000000000000001000";
  	pro(16) <= "00100000000010010000000000000101";
  	pro(17) <= "10101101000010010000000000000000";
  	pro(18) <= "00100001000010000000000000001000";
  	pro(19) <= "00100000000010010000000000000011";
  	pro(20) <= "10101101000010010000000000000000";
  	pro(21) <= "00100001000010000000000000001000";
  	pro(22) <= "00100000000010010000000000000001";
  	pro(23) <= "10101101000010010000000000000000";
  	pro(24) <= "00100001000010000000000000001000";
  	pro(25) <= "00100000000010010000000000000110";
  	pro(26) <= "10101101000010010000000000000000";
  	pro(27) <= "00100001000010000000000000001000";
  	pro(28) <= "00100000000010010000000000000000";
  	pro(29) <= "10101101000010010000000000000000";
  	pro(30) <= "00000000000000000100000000100000";
  	pro(31) <= "00100000000010010000000000101000";
  	pro(32) <= "00000001000010010111100000101010";
  	pro(33) <= "00010000000011110000000000001101";
  	pro(34) <= "00100001000010100000000000000100";
  	pro(35) <= "00000001010010010111100000101010";
  	pro(36) <= "00010000000011110000000000000111";
  	pro(37) <= "10001101000100000000000000000000";
  	pro(38) <= "10001101000100010000000000000000";
  	pro(39) <= "00000010001100000111100000101010";
  	pro(40) <= "00010000000011110000000000000010";
  	pro(41) <= "10101101000100010000000000000000";	
  	pro(42) <= "10101101010100000000000000000000";
  	pro(43) <= "00100001010010100000000000000100";
  	pro(44) <= "00001000000000000000000000100011";
  	pro(45) <= "00100001000010000000000000000100";
  	pro(46) <= "00001000000000000000000000100000";
  	pro(47) <= "00000000000000000000000000000000";
  	pro(48) <= "00000000000000000000000000000000";
  	pro(49) <= "00000000000000000000000000000000";
  	pro(50) <= "00000000000000000000000000000000";
  	pro(51) <= "00000000000000000000000000000000";
  	pro(52) <= "00000000000000000000000000000000";
  	pro(53) <= "00000000000000000000000000000000";
  	pro(54) <= "00000000000000000000000000000000";
  	pro(55) <= "00000000000000000000000000000000";
  	pro(56) <= "00000000000000000000000000000000";
  	pro(57) <= "00000000000000000000000000000000";
  	pro(58) <= "00000000000000000000000000000000";
  	pro(59) <= "00000000000000000000000000000000";
  	pro(60) <= "00000000000000000000000000000000";
  	pro(61) <= "00000000000000000000000000000000";
  	pro(62) <= "00000000000000000000000000000000";
  	pro(63) <= "00000000000000000000000000000000";
  	
  	for i in 0 to 10000 loop
  	  wait for 10 ns;
  	  clock <= '1';
  	  wait for 10 ns;
 	   clock <= '0';
   end loop;
  end process;
end cmp;
