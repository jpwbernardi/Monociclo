library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package NovosTipos is
  type VetorWord is array(natural range <>) of signed(31 downto 0);
end;
